package tartaruga_pkg;

///////////////////////////////////////////////////////////////////////////////
// TYPES
///////////////////////////////////////////////////////////////////////////////

    typedef logic [31:0] bus32_t;



endpackage

module dummy_imem 
import 
(
input bus32_t
)

package tartaruga_pkg;

///////////////////////////////////////////////////////////////////////////////
// PARAMETERS
///////////////////////////////////////////////////////////////////////////////

parameter IMEM_POS = 4096;


///////////////////////////////////////////////////////////////////////////////
// TYPES
///////////////////////////////////////////////////////////////////////////////

    typedef logic [31:0] bus32_t;



endpackage

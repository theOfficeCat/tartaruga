module decoder
    import tartaruga_pkg::*;
    import riscv_pkg::*;
(
    input bus32_t pc_i,
    input instruction_t instr_i,
    output instr_data_t instr_decoded_o
);

    //assign instr_decoded_o = '0;

    always_comb begin
        instr_decoded_o.pc = pc_i;
        instr_decoded_o.instr = instr_i;
        instr_decoded_o.addr_rs1 = instr_i.rtype.rs1;
        instr_decoded_o.addr_rs2 = instr_i.rtype.rs2;
        instr_decoded_o.addr_rd = instr_i.rtype.rd;
        
        case (instr_i.rtype.opcode)
            OP_ALU_I: begin
                instr_decoded_o.write_enable = 1'b1;
                instr_decoded_o.rs1_or_pc = RS1;
                instr_decoded_o.rs2_or_imm = IMM;
                instr_decoded_o.alu_or_mem = ALU;
                instr_decoded_o.store_to_mem = 1'b0;

                case (instr_i.rtype.func3)
                    F3_ADD_SUB: begin //ADDI
                        instr_decoded_o.alu_op = ADD;
                    end
                    F3_SLT: begin //SLTI
                        instr_decoded_o.alu_op = SLT;
                    end
                    F3_SLTU: begin //SLTIU
                        instr_decoded_o.alu_op = SLTU;
                    end
                    F3_XOR: begin //XORI
                        instr_decoded_o.alu_op = XOR;
                    end
                    F3_OR: begin //ORI
                        instr_decoded_o.alu_op = OR;
                    end
                    F3_AND: begin //ANDI
                        instr_decoded_o.alu_op = AND;
                    end
                    F3_SLL: begin //SLLI
                        case (instr_i.rtype.func7)
                            F7_ALU_NORMAL: begin
                                instr_decoded_o.alu_op = SLL;
                            end
                            default: begin
                                // illegal instruction treated as NOP being a x0 + x0
                                // without write

                                instr_decoded_o.write_enable = 1'b0;
                                instr_decoded_o.rs1_or_pc = RS1;
                                instr_decoded_o.rs2_or_imm = RS2;
                                instr_decoded_o.addr_rs1 = '0;
                                instr_decoded_o.addr_rs2 = '0;
                                instr_decoded_o.addr_rd = '0;
                                instr_decoded_o.alu_op = ADD;
                                instr_decoded_o.alu_or_mem = ALU;
                                instr_decoded_o.store_to_mem = 1'b0;
                            end
                        endcase
                    end
                    F3_SRL_SRA: begin //SRLI and SRAI
                        case (instr_i.rtype.func7)
                            F7_ALU_NORMAL: begin
                                instr_decoded_o.alu_op = SRL;
                            end
                            F7_ALU_MODIFIED: begin
                                instr_decoded_o.alu_op = SRA;
                            end
                            default: begin
                                // illegal instruction treated as NOP being a x0 + x0
                                // without write

                                instr_decoded_o.write_enable = 1'b0;
                                instr_decoded_o.rs1_or_pc = RS1;
                                instr_decoded_o.rs2_or_imm = RS2;
                                instr_decoded_o.addr_rs1 = '0;
                                instr_decoded_o.addr_rs2 = '0;
                                instr_decoded_o.addr_rd = '0;
                                instr_decoded_o.alu_op = ADD;
                                instr_decoded_o.alu_or_mem = ALU;
                                instr_decoded_o.store_to_mem = 1'b0;
                            end
                        endcase
                    end
                    default: begin
                        // illegal instruction treated as NOP being a x0 + x0
                        // without write

                        instr_decoded_o.write_enable = 1'b0;
                        instr_decoded_o.rs1_or_pc = RS1;
                        instr_decoded_o.rs2_or_imm = RS2;
                        instr_decoded_o.addr_rs1 = '0;
                        instr_decoded_o.addr_rs2 = '0;
                        instr_decoded_o.addr_rd = '0;
                        instr_decoded_o.alu_op = ADD;
                        instr_decoded_o.alu_or_mem = ALU;
                        instr_decoded_o.store_to_mem = 1'b0;
                    end
                endcase
            end

            OP_ALU: begin
                instr_decoded_o.write_enable = 1'b1;
                instr_decoded_o.rs1_or_pc = RS1;
                instr_decoded_o.rs2_or_imm = RS2;
                instr_decoded_o.alu_or_mem = ALU;
                instr_decoded_o.store_to_mem = 1'b0;

                case (instr_i.rtype.func3)
                    F3_ADD_SUB: begin
                        case (instr_i.rtype.func7)
                            F7_ALU_NORMAL: begin
                                instr_decoded_o.alu_op = ADD;
                            end
                            F7_ALU_MODIFIED: begin
                                instr_decoded_o.alu_op = SUB;
                            end
                            default: begin
                                // illegal instruction treated as NOP being a x0 + x0
                                // without write

                                instr_decoded_o.write_enable = 1'b0;
                                instr_decoded_o.rs1_or_pc = RS1;
                                instr_decoded_o.rs2_or_imm = RS2;
                                instr_decoded_o.addr_rs1 = '0;
                                instr_decoded_o.addr_rs2 = '0;
                                instr_decoded_o.addr_rd = '0;
                                instr_decoded_o.alu_op = ADD;
                                instr_decoded_o.alu_or_mem = ALU;
                                instr_decoded_o.store_to_mem = 1'b0;
                            end
                        endcase
                    end
                    F3_SLL: begin
                         case (instr_i.rtype.func7)
                            F7_ALU_NORMAL: begin
                                instr_decoded_o.alu_op = SLL;
                            end
                            default: begin
                                // illegal instruction treated as NOP being a x0 + x0
                                // without write

                                instr_decoded_o.write_enable = 1'b0;
                                instr_decoded_o.rs1_or_pc = RS1;
                                instr_decoded_o.rs2_or_imm = RS2;
                                instr_decoded_o.addr_rs1 = '0;
                                instr_decoded_o.addr_rs2 = '0;
                                instr_decoded_o.addr_rd = '0;
                                instr_decoded_o.alu_op = ADD;
                                instr_decoded_o.alu_or_mem = ALU;
                                instr_decoded_o.store_to_mem = 1'b0;
                            end
                        endcase
                    end
                    F3_SLT: begin
                         case (instr_i.rtype.func7)
                            F7_ALU_NORMAL: begin
                                instr_decoded_o.alu_op = SLT;
                            end
                            default: begin
                                // illegal instruction treated as NOP being a x0 + x0
                                // without write

                                instr_decoded_o.write_enable = 1'b0;
                                instr_decoded_o.rs1_or_pc = RS1;
                                instr_decoded_o.rs2_or_imm = RS2;
                                instr_decoded_o.addr_rs1 = '0;
                                instr_decoded_o.addr_rs2 = '0;
                                instr_decoded_o.addr_rd = '0;
                                instr_decoded_o.alu_op = ADD;
                                instr_decoded_o.alu_or_mem = ALU;
                                instr_decoded_o.store_to_mem = 1'b0;
                            end
                        endcase
                    end
                    F3_SLTU: begin
                         case (instr_i.rtype.func7)
                            F7_ALU_NORMAL: begin
                                instr_decoded_o.alu_op = SLTU;
                            end
                            default: begin
                                // illegal instruction treated as NOP being a x0 + x0
                                // without write

                                instr_decoded_o.write_enable = 1'b0;
                                instr_decoded_o.rs1_or_pc = RS1;
                                instr_decoded_o.rs2_or_imm = RS2;
                                instr_decoded_o.addr_rs1 = '0;
                                instr_decoded_o.addr_rs2 = '0;
                                instr_decoded_o.addr_rd = '0;
                                instr_decoded_o.alu_op = ADD;
                                instr_decoded_o.alu_or_mem = ALU;
                                instr_decoded_o.store_to_mem = 1'b0;
                            end
                        endcase
                    end
                    F3_XOR: begin
                         case (instr_i.rtype.func7)
                            F7_ALU_NORMAL: begin
                                instr_decoded_o.alu_op = XOR;
                            end
                            default: begin
                                // illegal instruction treated as NOP being a x0 + x0
                                // without write

                                instr_decoded_o.write_enable = 1'b0;
                                instr_decoded_o.rs1_or_pc = RS1;
                                instr_decoded_o.rs2_or_imm = RS2;
                                instr_decoded_o.addr_rs1 = '0;
                                instr_decoded_o.addr_rs2 = '0;
                                instr_decoded_o.addr_rd = '0;
                                instr_decoded_o.alu_op = ADD;
                                instr_decoded_o.alu_or_mem = ALU;
                                instr_decoded_o.store_to_mem = 1'b0;
                            end
                        endcase
                    end
                    F3_SRL_SRA: begin
                         case (instr_i.rtype.func7)
                            F7_ALU_NORMAL: begin
                                instr_decoded_o.alu_op = SRL;
                            end
                            F7_ALU_MODIFIED: begin
                                instr_decoded_o.alu_op = SRA;
                            end
                            default: begin
                                // illegal instruction treated as NOP being a x0 + x0
                                // without write

                                instr_decoded_o.write_enable = 1'b0;
                                instr_decoded_o.rs1_or_pc = RS1;
                                instr_decoded_o.rs2_or_imm = RS2;
                                instr_decoded_o.addr_rs1 = '0;
                                instr_decoded_o.addr_rs2 = '0;
                                instr_decoded_o.addr_rd = '0;
                                instr_decoded_o.alu_op = ADD;
                                instr_decoded_o.alu_or_mem = ALU;
                                instr_decoded_o.store_to_mem = 1'b0;
                            end
                        endcase
                    end
                    F3_OR: begin
                         case (instr_i.rtype.func7)
                            F7_ALU_NORMAL: begin
                                instr_decoded_o.alu_op = OR;
                            end
                            default: begin
                                // illegal instruction treated as NOP being a x0 + x0
                                // without write

                                instr_decoded_o.write_enable = 1'b0;
                                instr_decoded_o.rs1_or_pc = RS1;
                                instr_decoded_o.rs2_or_imm = RS2;
                                instr_decoded_o.addr_rs1 = '0;
                                instr_decoded_o.addr_rs2 = '0;
                                instr_decoded_o.addr_rd = '0;
                                instr_decoded_o.alu_op = ADD;
                                instr_decoded_o.alu_or_mem = ALU;
                                instr_decoded_o.store_to_mem = 1'b0;
                            end
                        endcase
                    end
                    F3_AND: begin
                         case (instr_i.rtype.func7)
                            F7_ALU_NORMAL: begin
                                instr_decoded_o.alu_op = AND;
                            end
                            default: begin
                                // illegal instruction treated as NOP being a x0 + x0
                                // without write

                                instr_decoded_o.write_enable = 1'b0;
                                instr_decoded_o.rs1_or_pc = RS1;
                                instr_decoded_o.rs2_or_imm = RS2;
                                instr_decoded_o.addr_rs1 = '0;
                                instr_decoded_o.addr_rs2 = '0;
                                instr_decoded_o.addr_rd = '0;
                                instr_decoded_o.alu_op = ADD;
                                instr_decoded_o.alu_or_mem = ALU;
                                instr_decoded_o.store_to_mem = 1'b0;
                            end
                        endcase
                    end
 
                    default: begin
                        // illegal instruction treated as NOP being a x0 + x0
                        // without write

                        instr_decoded_o.write_enable = 1'b0;
                        instr_decoded_o.rs1_or_pc = RS1;
                        instr_decoded_o.rs2_or_imm = RS2;
                        instr_decoded_o.addr_rs1 = '0;
                        instr_decoded_o.addr_rs2 = '0;
                        instr_decoded_o.addr_rd = '0;
                        instr_decoded_o.alu_op = ADD;
                        instr_decoded_o.store_to_mem = 1'b0;
                    end
                endcase
            end

            OP_LUI: begin
                instr_decoded_o.write_enable = 1'b1;
                instr_decoded_o.rs1_or_pc = RS1;
                instr_decoded_o.rs2_or_imm = IMM;
                instr_decoded_o.alu_op = ADD;
                instr_decoded_o.alu_or_mem = ALU;
                instr_decoded_o.store_to_mem = 1'b0;

                instr_decoded_o.addr_rs1 = '0; // Hardcoded to x0 which is hardwired to 0
            end

            OP_AUIPC: begin
                instr_decoded_o.write_enable = 1'b1;
                instr_decoded_o.rs1_or_pc = PC;
                instr_decoded_o.rs2_or_imm = IMM;
                instr_decoded_o.alu_op = ADD;
                instr_decoded_o.alu_or_mem = ALU;
                instr_decoded_o.store_to_mem = 1'b0;
            end
            default: begin
                // illegal instruction treated as NOP being a x0 + x0
                // without write

                instr_decoded_o.write_enable = 1'b0;
                instr_decoded_o.rs1_or_pc = RS1;
                instr_decoded_o.rs2_or_imm = RS2;
                instr_decoded_o.addr_rs1 = '0;
                instr_decoded_o.addr_rs2 = '0;
                instr_decoded_o.addr_rd = '0;
                instr_decoded_o.alu_op = ADD;
                instr_decoded_o.alu_or_mem = ALU;
                instr_decoded_o.store_to_mem = 1'b0;
            end
        endcase
    end

endmodule

module scoreboard
    import tartaruga_pkg::*;
(
    
);

// Input decode_to_exe enters on number of cycles on exe - 1:
// - Index 3 on multiplications
// - Index 0 on the other ones
//
// Unit releases index 0
// If instruction on the index is already valid stall decode and fetch this
// cycle

endmodule

module top
(

);


endmodule
